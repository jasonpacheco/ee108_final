module sine_rom (
    input clk,
    input [9:0] addr,
    output reg [15:0] dout
);

    wire [15:0] memory [1023:0];

    always @(posedge clk)
        dout = memory[addr];

    assign memory[    0 ] = 16'd00000;
    assign memory[    1 ] = 16'd00050;
    assign memory[    2 ] = 16'd00101;
    assign memory[    3 ] = 16'd00151;
    assign memory[    4 ] = 16'd00201;
    assign memory[    5 ] = 16'd00251;
    assign memory[    6 ] = 16'd00302;
    assign memory[    7 ] = 16'd00352;
    assign memory[    8 ] = 16'd00402;
    assign memory[    9 ] = 16'd00452;
    assign memory[   10 ] = 16'd00503;
    assign memory[   11 ] = 16'd00553;
    assign memory[   12 ] = 16'd00603;
    assign memory[   13 ] = 16'd00653;
    assign memory[   14 ] = 16'd00704;
    assign memory[   15 ] = 16'd00754;
    assign memory[   16 ] = 16'd00804;
    assign memory[   17 ] = 16'd00854;
    assign memory[   18 ] = 16'd00905;
    assign memory[   19 ] = 16'd00955;
    assign memory[   20 ] = 16'd01005;
    assign memory[   21 ] = 16'd01055;
    assign memory[   22 ] = 16'd01106;
    assign memory[   23 ] = 16'd01156;
    assign memory[   24 ] = 16'd01206;
    assign memory[   25 ] = 16'd01256;
    assign memory[   26 ] = 16'd01307;
    assign memory[   27 ] = 16'd01357;
    assign memory[   28 ] = 16'd01407;
    assign memory[   29 ] = 16'd01457;
    assign memory[   30 ] = 16'd01507;
    assign memory[   31 ] = 16'd01558;
    assign memory[   32 ] = 16'd01608;
    assign memory[   33 ] = 16'd01658;
    assign memory[   34 ] = 16'd01708;
    assign memory[   35 ] = 16'd01758;
    assign memory[   36 ] = 16'd01809;
    assign memory[   37 ] = 16'd01859;
    assign memory[   38 ] = 16'd01909;
    assign memory[   39 ] = 16'd01959;
    assign memory[   40 ] = 16'd02009;
    assign memory[   41 ] = 16'd02059;
    assign memory[   42 ] = 16'd02110;
    assign memory[   43 ] = 16'd02160;
    assign memory[   44 ] = 16'd02210;
    assign memory[   45 ] = 16'd02260;
    assign memory[   46 ] = 16'd02310;
    assign memory[   47 ] = 16'd02360;
    assign memory[   48 ] = 16'd02410;
    assign memory[   49 ] = 16'd02461;
    assign memory[   50 ] = 16'd02511;
    assign memory[   51 ] = 16'd02561;
    assign memory[   52 ] = 16'd02611;
    assign memory[   53 ] = 16'd02661;
    assign memory[   54 ] = 16'd02711;
    assign memory[   55 ] = 16'd02761;
    assign memory[   56 ] = 16'd02811;
    assign memory[   57 ] = 16'd02861;
    assign memory[   58 ] = 16'd02911;
    assign memory[   59 ] = 16'd02962;
    assign memory[   60 ] = 16'd03012;
    assign memory[   61 ] = 16'd03062;
    assign memory[   62 ] = 16'd03112;
    assign memory[   63 ] = 16'd03162;
    assign memory[   64 ] = 16'd03212;
    assign memory[   65 ] = 16'd03262;
    assign memory[   66 ] = 16'd03312;
    assign memory[   67 ] = 16'd03362;
    assign memory[   68 ] = 16'd03412;
    assign memory[   69 ] = 16'd03462;
    assign memory[   70 ] = 16'd03512;
    assign memory[   71 ] = 16'd03562;
    assign memory[   72 ] = 16'd03612;
    assign memory[   73 ] = 16'd03662;
    assign memory[   74 ] = 16'd03712;
    assign memory[   75 ] = 16'd03761;
    assign memory[   76 ] = 16'd03811;
    assign memory[   77 ] = 16'd03861;
    assign memory[   78 ] = 16'd03911;
    assign memory[   79 ] = 16'd03961;
    assign memory[   80 ] = 16'd04011;
    assign memory[   81 ] = 16'd04061;
    assign memory[   82 ] = 16'd04111;
    assign memory[   83 ] = 16'd04161;
    assign memory[   84 ] = 16'd04210;
    assign memory[   85 ] = 16'd04260;
    assign memory[   86 ] = 16'd04310;
    assign memory[   87 ] = 16'd04360;
    assign memory[   88 ] = 16'd04410;
    assign memory[   89 ] = 16'd04460;
    assign memory[   90 ] = 16'd04509;
    assign memory[   91 ] = 16'd04559;
    assign memory[   92 ] = 16'd04609;
    assign memory[   93 ] = 16'd04659;
    assign memory[   94 ] = 16'd04708;
    assign memory[   95 ] = 16'd04758;
    assign memory[   96 ] = 16'd04808;
    assign memory[   97 ] = 16'd04858;
    assign memory[   98 ] = 16'd04907;
    assign memory[   99 ] = 16'd04957;
    assign memory[  100 ] = 16'd05007;
    assign memory[  101 ] = 16'd05056;
    assign memory[  102 ] = 16'd05106;
    assign memory[  103 ] = 16'd05156;
    assign memory[  104 ] = 16'd05205;
    assign memory[  105 ] = 16'd05255;
    assign memory[  106 ] = 16'd05305;
    assign memory[  107 ] = 16'd05354;
    assign memory[  108 ] = 16'd05404;
    assign memory[  109 ] = 16'd05453;
    assign memory[  110 ] = 16'd05503;
    assign memory[  111 ] = 16'd05552;
    assign memory[  112 ] = 16'd05602;
    assign memory[  113 ] = 16'd05651;
    assign memory[  114 ] = 16'd05701;
    assign memory[  115 ] = 16'd05750;
    assign memory[  116 ] = 16'd05800;
    assign memory[  117 ] = 16'd05849;
    assign memory[  118 ] = 16'd05899;
    assign memory[  119 ] = 16'd05948;
    assign memory[  120 ] = 16'd05998;
    assign memory[  121 ] = 16'd06047;
    assign memory[  122 ] = 16'd06096;
    assign memory[  123 ] = 16'd06146;
    assign memory[  124 ] = 16'd06195;
    assign memory[  125 ] = 16'd06245;
    assign memory[  126 ] = 16'd06294;
    assign memory[  127 ] = 16'd06343;
    assign memory[  128 ] = 16'd06393;
    assign memory[  129 ] = 16'd06442;
    assign memory[  130 ] = 16'd06491;
    assign memory[  131 ] = 16'd06540;
    assign memory[  132 ] = 16'd06590;
    assign memory[  133 ] = 16'd06639;
    assign memory[  134 ] = 16'd06688;
    assign memory[  135 ] = 16'd06737;
    assign memory[  136 ] = 16'd06786;
    assign memory[  137 ] = 16'd06836;
    assign memory[  138 ] = 16'd06885;
    assign memory[  139 ] = 16'd06934;
    assign memory[  140 ] = 16'd06983;
    assign memory[  141 ] = 16'd07032;
    assign memory[  142 ] = 16'd07081;
    assign memory[  143 ] = 16'd07130;
    assign memory[  144 ] = 16'd07179;
    assign memory[  145 ] = 16'd07228;
    assign memory[  146 ] = 16'd07277;
    assign memory[  147 ] = 16'd07326;
    assign memory[  148 ] = 16'd07375;
    assign memory[  149 ] = 16'd07424;
    assign memory[  150 ] = 16'd07473;
    assign memory[  151 ] = 16'd07522;
    assign memory[  152 ] = 16'd07571;
    assign memory[  153 ] = 16'd07620;
    assign memory[  154 ] = 16'd07669;
    assign memory[  155 ] = 16'd07718;
    assign memory[  156 ] = 16'd07767;
    assign memory[  157 ] = 16'd07815;
    assign memory[  158 ] = 16'd07864;
    assign memory[  159 ] = 16'd07913;
    assign memory[  160 ] = 16'd07962;
    assign memory[  161 ] = 16'd08010;
    assign memory[  162 ] = 16'd08059;
    assign memory[  163 ] = 16'd08108;
    assign memory[  164 ] = 16'd08157;
    assign memory[  165 ] = 16'd08205;
    assign memory[  166 ] = 16'd08254;
    assign memory[  167 ] = 16'd08303;
    assign memory[  168 ] = 16'd08351;
    assign memory[  169 ] = 16'd08400;
    assign memory[  170 ] = 16'd08448;
    assign memory[  171 ] = 16'd08497;
    assign memory[  172 ] = 16'd08545;
    assign memory[  173 ] = 16'd08594;
    assign memory[  174 ] = 16'd08642;
    assign memory[  175 ] = 16'd08691;
    assign memory[  176 ] = 16'd08739;
    assign memory[  177 ] = 16'd08788;
    assign memory[  178 ] = 16'd08836;
    assign memory[  179 ] = 16'd08885;
    assign memory[  180 ] = 16'd08933;
    assign memory[  181 ] = 16'd08981;
    assign memory[  182 ] = 16'd09030;
    assign memory[  183 ] = 16'd09078;
    assign memory[  184 ] = 16'd09126;
    assign memory[  185 ] = 16'd09175;
    assign memory[  186 ] = 16'd09223;
    assign memory[  187 ] = 16'd09271;
    assign memory[  188 ] = 16'd09319;
    assign memory[  189 ] = 16'd09367;
    assign memory[  190 ] = 16'd09416;
    assign memory[  191 ] = 16'd09464;
    assign memory[  192 ] = 16'd09512;
    assign memory[  193 ] = 16'd09560;
    assign memory[  194 ] = 16'd09608;
    assign memory[  195 ] = 16'd09656;
    assign memory[  196 ] = 16'd09704;
    assign memory[  197 ] = 16'd09752;
    assign memory[  198 ] = 16'd09800;
    assign memory[  199 ] = 16'd09848;
    assign memory[  200 ] = 16'd09896;
    assign memory[  201 ] = 16'd09944;
    assign memory[  202 ] = 16'd09992;
    assign memory[  203 ] = 16'd10039;
    assign memory[  204 ] = 16'd10087;
    assign memory[  205 ] = 16'd10135;
    assign memory[  206 ] = 16'd10183;
    assign memory[  207 ] = 16'd10231;
    assign memory[  208 ] = 16'd10278;
    assign memory[  209 ] = 16'd10326;
    assign memory[  210 ] = 16'd10374;
    assign memory[  211 ] = 16'd10421;
    assign memory[  212 ] = 16'd10469;
    assign memory[  213 ] = 16'd10517;
    assign memory[  214 ] = 16'd10564;
    assign memory[  215 ] = 16'd10612;
    assign memory[  216 ] = 16'd10659;
    assign memory[  217 ] = 16'd10707;
    assign memory[  218 ] = 16'd10754;
    assign memory[  219 ] = 16'd10802;
    assign memory[  220 ] = 16'd10849;
    assign memory[  221 ] = 16'd10897;
    assign memory[  222 ] = 16'd10944;
    assign memory[  223 ] = 16'd10992;
    assign memory[  224 ] = 16'd11039;
    assign memory[  225 ] = 16'd11086;
    assign memory[  226 ] = 16'd11133;
    assign memory[  227 ] = 16'd11181;
    assign memory[  228 ] = 16'd11228;
    assign memory[  229 ] = 16'd11275;
    assign memory[  230 ] = 16'd11322;
    assign memory[  231 ] = 16'd11370;
    assign memory[  232 ] = 16'd11417;
    assign memory[  233 ] = 16'd11464;
    assign memory[  234 ] = 16'd11511;
    assign memory[  235 ] = 16'd11558;
    assign memory[  236 ] = 16'd11605;
    assign memory[  237 ] = 16'd11652;
    assign memory[  238 ] = 16'd11699;
    assign memory[  239 ] = 16'd11746;
    assign memory[  240 ] = 16'd11793;
    assign memory[  241 ] = 16'd11840;
    assign memory[  242 ] = 16'd11886;
    assign memory[  243 ] = 16'd11933;
    assign memory[  244 ] = 16'd11980;
    assign memory[  245 ] = 16'd12027;
    assign memory[  246 ] = 16'd12074;
    assign memory[  247 ] = 16'd12120;
    assign memory[  248 ] = 16'd12167;
    assign memory[  249 ] = 16'd12214;
    assign memory[  250 ] = 16'd12260;
    assign memory[  251 ] = 16'd12307;
    assign memory[  252 ] = 16'd12353;
    assign memory[  253 ] = 16'd12400;
    assign memory[  254 ] = 16'd12446;
    assign memory[  255 ] = 16'd12493;
    assign memory[  256 ] = 16'd12539;
    assign memory[  257 ] = 16'd12586;
    assign memory[  258 ] = 16'd12632;
    assign memory[  259 ] = 16'd12679;
    assign memory[  260 ] = 16'd12725;
    assign memory[  261 ] = 16'd12771;
    assign memory[  262 ] = 16'd12817;
    assign memory[  263 ] = 16'd12864;
    assign memory[  264 ] = 16'd12910;
    assign memory[  265 ] = 16'd12956;
    assign memory[  266 ] = 16'd13002;
    assign memory[  267 ] = 16'd13048;
    assign memory[  268 ] = 16'd13094;
    assign memory[  269 ] = 16'd13141;
    assign memory[  270 ] = 16'd13187;
    assign memory[  271 ] = 16'd13233;
    assign memory[  272 ] = 16'd13279;
    assign memory[  273 ] = 16'd13324;
    assign memory[  274 ] = 16'd13370;
    assign memory[  275 ] = 16'd13416;
    assign memory[  276 ] = 16'd13462;
    assign memory[  277 ] = 16'd13508;
    assign memory[  278 ] = 16'd13554;
    assign memory[  279 ] = 16'd13599;
    assign memory[  280 ] = 16'd13645;
    assign memory[  281 ] = 16'd13691;
    assign memory[  282 ] = 16'd13736;
    assign memory[  283 ] = 16'd13782;
    assign memory[  284 ] = 16'd13828;
    assign memory[  285 ] = 16'd13873;
    assign memory[  286 ] = 16'd13919;
    assign memory[  287 ] = 16'd13964;
    assign memory[  288 ] = 16'd14010;
    assign memory[  289 ] = 16'd14055;
    assign memory[  290 ] = 16'd14101;
    assign memory[  291 ] = 16'd14146;
    assign memory[  292 ] = 16'd14191;
    assign memory[  293 ] = 16'd14236;
    assign memory[  294 ] = 16'd14282;
    assign memory[  295 ] = 16'd14327;
    assign memory[  296 ] = 16'd14372;
    assign memory[  297 ] = 16'd14417;
    assign memory[  298 ] = 16'd14462;
    assign memory[  299 ] = 16'd14507;
    assign memory[  300 ] = 16'd14553;
    assign memory[  301 ] = 16'd14598;
    assign memory[  302 ] = 16'd14643;
    assign memory[  303 ] = 16'd14688;
    assign memory[  304 ] = 16'd14732;
    assign memory[  305 ] = 16'd14777;
    assign memory[  306 ] = 16'd14822;
    assign memory[  307 ] = 16'd14867;
    assign memory[  308 ] = 16'd14912;
    assign memory[  309 ] = 16'd14956;
    assign memory[  310 ] = 16'd15001;
    assign memory[  311 ] = 16'd15046;
    assign memory[  312 ] = 16'd15090;
    assign memory[  313 ] = 16'd15135;
    assign memory[  314 ] = 16'd15180;
    assign memory[  315 ] = 16'd15224;
    assign memory[  316 ] = 16'd15269;
    assign memory[  317 ] = 16'd15313;
    assign memory[  318 ] = 16'd15358;
    assign memory[  319 ] = 16'd15402;
    assign memory[  320 ] = 16'd15446;
    assign memory[  321 ] = 16'd15491;
    assign memory[  322 ] = 16'd15535;
    assign memory[  323 ] = 16'd15579;
    assign memory[  324 ] = 16'd15623;
    assign memory[  325 ] = 16'd15667;
    assign memory[  326 ] = 16'd15712;
    assign memory[  327 ] = 16'd15756;
    assign memory[  328 ] = 16'd15800;
    assign memory[  329 ] = 16'd15844;
    assign memory[  330 ] = 16'd15888;
    assign memory[  331 ] = 16'd15932;
    assign memory[  332 ] = 16'd15976;
    assign memory[  333 ] = 16'd16019;
    assign memory[  334 ] = 16'd16063;
    assign memory[  335 ] = 16'd16107;
    assign memory[  336 ] = 16'd16151;
    assign memory[  337 ] = 16'd16195;
    assign memory[  338 ] = 16'd16238;
    assign memory[  339 ] = 16'd16282;
    assign memory[  340 ] = 16'd16325;
    assign memory[  341 ] = 16'd16369;
    assign memory[  342 ] = 16'd16413;
    assign memory[  343 ] = 16'd16456;
    assign memory[  344 ] = 16'd16499;
    assign memory[  345 ] = 16'd16543;
    assign memory[  346 ] = 16'd16586;
    assign memory[  347 ] = 16'd16630;
    assign memory[  348 ] = 16'd16673;
    assign memory[  349 ] = 16'd16716;
    assign memory[  350 ] = 16'd16759;
    assign memory[  351 ] = 16'd16802;
    assign memory[  352 ] = 16'd16846;
    assign memory[  353 ] = 16'd16889;
    assign memory[  354 ] = 16'd16932;
    assign memory[  355 ] = 16'd16975;
    assign memory[  356 ] = 16'd17018;
    assign memory[  357 ] = 16'd17061;
    assign memory[  358 ] = 16'd17104;
    assign memory[  359 ] = 16'd17146;
    assign memory[  360 ] = 16'd17189;
    assign memory[  361 ] = 16'd17232;
    assign memory[  362 ] = 16'd17275;
    assign memory[  363 ] = 16'd17317;
    assign memory[  364 ] = 16'd17360;
    assign memory[  365 ] = 16'd17403;
    assign memory[  366 ] = 16'd17445;
    assign memory[  367 ] = 16'd17488;
    assign memory[  368 ] = 16'd17530;
    assign memory[  369 ] = 16'd17573;
    assign memory[  370 ] = 16'd17615;
    assign memory[  371 ] = 16'd17657;
    assign memory[  372 ] = 16'd17700;
    assign memory[  373 ] = 16'd17742;
    assign memory[  374 ] = 16'd17784;
    assign memory[  375 ] = 16'd17827;
    assign memory[  376 ] = 16'd17869;
    assign memory[  377 ] = 16'd17911;
    assign memory[  378 ] = 16'd17953;
    assign memory[  379 ] = 16'd17995;
    assign memory[  380 ] = 16'd18037;
    assign memory[  381 ] = 16'd18079;
    assign memory[  382 ] = 16'd18121;
    assign memory[  383 ] = 16'd18163;
    assign memory[  384 ] = 16'd18204;
    assign memory[  385 ] = 16'd18246;
    assign memory[  386 ] = 16'd18288;
    assign memory[  387 ] = 16'd18330;
    assign memory[  388 ] = 16'd18371;
    assign memory[  389 ] = 16'd18413;
    assign memory[  390 ] = 16'd18454;
    assign memory[  391 ] = 16'd18496;
    assign memory[  392 ] = 16'd18537;
    assign memory[  393 ] = 16'd18579;
    assign memory[  394 ] = 16'd18620;
    assign memory[  395 ] = 16'd18661;
    assign memory[  396 ] = 16'd18703;
    assign memory[  397 ] = 16'd18744;
    assign memory[  398 ] = 16'd18785;
    assign memory[  399 ] = 16'd18826;
    assign memory[  400 ] = 16'd18868;
    assign memory[  401 ] = 16'd18909;
    assign memory[  402 ] = 16'd18950;
    assign memory[  403 ] = 16'd18991;
    assign memory[  404 ] = 16'd19032;
    assign memory[  405 ] = 16'd19072;
    assign memory[  406 ] = 16'd19113;
    assign memory[  407 ] = 16'd19154;
    assign memory[  408 ] = 16'd19195;
    assign memory[  409 ] = 16'd19236;
    assign memory[  410 ] = 16'd19276;
    assign memory[  411 ] = 16'd19317;
    assign memory[  412 ] = 16'd19357;
    assign memory[  413 ] = 16'd19398;
    assign memory[  414 ] = 16'd19438;
    assign memory[  415 ] = 16'd19479;
    assign memory[  416 ] = 16'd19519;
    assign memory[  417 ] = 16'd19560;
    assign memory[  418 ] = 16'd19600;
    assign memory[  419 ] = 16'd19640;
    assign memory[  420 ] = 16'd19680;
    assign memory[  421 ] = 16'd19721;
    assign memory[  422 ] = 16'd19761;
    assign memory[  423 ] = 16'd19801;
    assign memory[  424 ] = 16'd19841;
    assign memory[  425 ] = 16'd19881;
    assign memory[  426 ] = 16'd19921;
    assign memory[  427 ] = 16'd19961;
    assign memory[  428 ] = 16'd20000;
    assign memory[  429 ] = 16'd20040;
    assign memory[  430 ] = 16'd20080;
    assign memory[  431 ] = 16'd20120;
    assign memory[  432 ] = 16'd20159;
    assign memory[  433 ] = 16'd20199;
    assign memory[  434 ] = 16'd20238;
    assign memory[  435 ] = 16'd20278;
    assign memory[  436 ] = 16'd20317;
    assign memory[  437 ] = 16'd20357;
    assign memory[  438 ] = 16'd20396;
    assign memory[  439 ] = 16'd20436;
    assign memory[  440 ] = 16'd20475;
    assign memory[  441 ] = 16'd20514;
    assign memory[  442 ] = 16'd20553;
    assign memory[  443 ] = 16'd20592;
    assign memory[  444 ] = 16'd20631;
    assign memory[  445 ] = 16'd20670;
    assign memory[  446 ] = 16'd20709;
    assign memory[  447 ] = 16'd20748;
    assign memory[  448 ] = 16'd20787;
    assign memory[  449 ] = 16'd20826;
    assign memory[  450 ] = 16'd20865;
    assign memory[  451 ] = 16'd20904;
    assign memory[  452 ] = 16'd20942;
    assign memory[  453 ] = 16'd20981;
    assign memory[  454 ] = 16'd21019;
    assign memory[  455 ] = 16'd21058;
    assign memory[  456 ] = 16'd21096;
    assign memory[  457 ] = 16'd21135;
    assign memory[  458 ] = 16'd21173;
    assign memory[  459 ] = 16'd21212;
    assign memory[  460 ] = 16'd21250;
    assign memory[  461 ] = 16'd21288;
    assign memory[  462 ] = 16'd21326;
    assign memory[  463 ] = 16'd21364;
    assign memory[  464 ] = 16'd21403;
    assign memory[  465 ] = 16'd21441;
    assign memory[  466 ] = 16'd21479;
    assign memory[  467 ] = 16'd21516;
    assign memory[  468 ] = 16'd21554;
    assign memory[  469 ] = 16'd21592;
    assign memory[  470 ] = 16'd21630;
    assign memory[  471 ] = 16'd21668;
    assign memory[  472 ] = 16'd21705;
    assign memory[  473 ] = 16'd21743;
    assign memory[  474 ] = 16'd21781;
    assign memory[  475 ] = 16'd21818;
    assign memory[  476 ] = 16'd21856;
    assign memory[  477 ] = 16'd21893;
    assign memory[  478 ] = 16'd21930;
    assign memory[  479 ] = 16'd21968;
    assign memory[  480 ] = 16'd22005;
    assign memory[  481 ] = 16'd22042;
    assign memory[  482 ] = 16'd22079;
    assign memory[  483 ] = 16'd22116;
    assign memory[  484 ] = 16'd22154;
    assign memory[  485 ] = 16'd22191;
    assign memory[  486 ] = 16'd22227;
    assign memory[  487 ] = 16'd22264;
    assign memory[  488 ] = 16'd22301;
    assign memory[  489 ] = 16'd22338;
    assign memory[  490 ] = 16'd22375;
    assign memory[  491 ] = 16'd22411;
    assign memory[  492 ] = 16'd22448;
    assign memory[  493 ] = 16'd22485;
    assign memory[  494 ] = 16'd22521;
    assign memory[  495 ] = 16'd22558;
    assign memory[  496 ] = 16'd22594;
    assign memory[  497 ] = 16'd22631;
    assign memory[  498 ] = 16'd22667;
    assign memory[  499 ] = 16'd22703;
    assign memory[  500 ] = 16'd22739;
    assign memory[  501 ] = 16'd22776;
    assign memory[  502 ] = 16'd22812;
    assign memory[  503 ] = 16'd22848;
    assign memory[  504 ] = 16'd22884;
    assign memory[  505 ] = 16'd22920;
    assign memory[  506 ] = 16'd22956;
    assign memory[  507 ] = 16'd22991;
    assign memory[  508 ] = 16'd23027;
    assign memory[  509 ] = 16'd23063;
    assign memory[  510 ] = 16'd23099;
    assign memory[  511 ] = 16'd23134;
    assign memory[  512 ] = 16'd23170;
    assign memory[  513 ] = 16'd23205;
    assign memory[  514 ] = 16'd23241;
    assign memory[  515 ] = 16'd23276;
    assign memory[  516 ] = 16'd23311;
    assign memory[  517 ] = 16'd23347;
    assign memory[  518 ] = 16'd23382;
    assign memory[  519 ] = 16'd23417;
    assign memory[  520 ] = 16'd23452;
    assign memory[  521 ] = 16'd23487;
    assign memory[  522 ] = 16'd23522;
    assign memory[  523 ] = 16'd23557;
    assign memory[  524 ] = 16'd23592;
    assign memory[  525 ] = 16'd23627;
    assign memory[  526 ] = 16'd23662;
    assign memory[  527 ] = 16'd23697;
    assign memory[  528 ] = 16'd23731;
    assign memory[  529 ] = 16'd23766;
    assign memory[  530 ] = 16'd23801;
    assign memory[  531 ] = 16'd23835;
    assign memory[  532 ] = 16'd23870;
    assign memory[  533 ] = 16'd23904;
    assign memory[  534 ] = 16'd23938;
    assign memory[  535 ] = 16'd23973;
    assign memory[  536 ] = 16'd24007;
    assign memory[  537 ] = 16'd24041;
    assign memory[  538 ] = 16'd24075;
    assign memory[  539 ] = 16'd24109;
    assign memory[  540 ] = 16'd24143;
    assign memory[  541 ] = 16'd24177;
    assign memory[  542 ] = 16'd24211;
    assign memory[  543 ] = 16'd24245;
    assign memory[  544 ] = 16'd24279;
    assign memory[  545 ] = 16'd24312;
    assign memory[  546 ] = 16'd24346;
    assign memory[  547 ] = 16'd24380;
    assign memory[  548 ] = 16'd24413;
    assign memory[  549 ] = 16'd24447;
    assign memory[  550 ] = 16'd24480;
    assign memory[  551 ] = 16'd24514;
    assign memory[  552 ] = 16'd24547;
    assign memory[  553 ] = 16'd24580;
    assign memory[  554 ] = 16'd24613;
    assign memory[  555 ] = 16'd24647;
    assign memory[  556 ] = 16'd24680;
    assign memory[  557 ] = 16'd24713;
    assign memory[  558 ] = 16'd24746;
    assign memory[  559 ] = 16'd24779;
    assign memory[  560 ] = 16'd24811;
    assign memory[  561 ] = 16'd24844;
    assign memory[  562 ] = 16'd24877;
    assign memory[  563 ] = 16'd24910;
    assign memory[  564 ] = 16'd24942;
    assign memory[  565 ] = 16'd24975;
    assign memory[  566 ] = 16'd25007;
    assign memory[  567 ] = 16'd25040;
    assign memory[  568 ] = 16'd25072;
    assign memory[  569 ] = 16'd25105;
    assign memory[  570 ] = 16'd25137;
    assign memory[  571 ] = 16'd25169;
    assign memory[  572 ] = 16'd25201;
    assign memory[  573 ] = 16'd25233;
    assign memory[  574 ] = 16'd25265;
    assign memory[  575 ] = 16'd25297;
    assign memory[  576 ] = 16'd25329;
    assign memory[  577 ] = 16'd25361;
    assign memory[  578 ] = 16'd25393;
    assign memory[  579 ] = 16'd25425;
    assign memory[  580 ] = 16'd25456;
    assign memory[  581 ] = 16'd25488;
    assign memory[  582 ] = 16'd25519;
    assign memory[  583 ] = 16'd25551;
    assign memory[  584 ] = 16'd25582;
    assign memory[  585 ] = 16'd25614;
    assign memory[  586 ] = 16'd25645;
    assign memory[  587 ] = 16'd25676;
    assign memory[  588 ] = 16'd25708;
    assign memory[  589 ] = 16'd25739;
    assign memory[  590 ] = 16'd25770;
    assign memory[  591 ] = 16'd25801;
    assign memory[  592 ] = 16'd25832;
    assign memory[  593 ] = 16'd25863;
    assign memory[  594 ] = 16'd25893;
    assign memory[  595 ] = 16'd25924;
    assign memory[  596 ] = 16'd25955;
    assign memory[  597 ] = 16'd25986;
    assign memory[  598 ] = 16'd26016;
    assign memory[  599 ] = 16'd26047;
    assign memory[  600 ] = 16'd26077;
    assign memory[  601 ] = 16'd26108;
    assign memory[  602 ] = 16'd26138;
    assign memory[  603 ] = 16'd26168;
    assign memory[  604 ] = 16'd26198;
    assign memory[  605 ] = 16'd26229;
    assign memory[  606 ] = 16'd26259;
    assign memory[  607 ] = 16'd26289;
    assign memory[  608 ] = 16'd26319;
    assign memory[  609 ] = 16'd26349;
    assign memory[  610 ] = 16'd26378;
    assign memory[  611 ] = 16'd26408;
    assign memory[  612 ] = 16'd26438;
    assign memory[  613 ] = 16'd26468;
    assign memory[  614 ] = 16'd26497;
    assign memory[  615 ] = 16'd26527;
    assign memory[  616 ] = 16'd26556;
    assign memory[  617 ] = 16'd26586;
    assign memory[  618 ] = 16'd26615;
    assign memory[  619 ] = 16'd26644;
    assign memory[  620 ] = 16'd26674;
    assign memory[  621 ] = 16'd26703;
    assign memory[  622 ] = 16'd26732;
    assign memory[  623 ] = 16'd26761;
    assign memory[  624 ] = 16'd26790;
    assign memory[  625 ] = 16'd26819;
    assign memory[  626 ] = 16'd26848;
    assign memory[  627 ] = 16'd26876;
    assign memory[  628 ] = 16'd26905;
    assign memory[  629 ] = 16'd26934;
    assign memory[  630 ] = 16'd26962;
    assign memory[  631 ] = 16'd26991;
    assign memory[  632 ] = 16'd27019;
    assign memory[  633 ] = 16'd27048;
    assign memory[  634 ] = 16'd27076;
    assign memory[  635 ] = 16'd27104;
    assign memory[  636 ] = 16'd27133;
    assign memory[  637 ] = 16'd27161;
    assign memory[  638 ] = 16'd27189;
    assign memory[  639 ] = 16'd27217;
    assign memory[  640 ] = 16'd27245;
    assign memory[  641 ] = 16'd27273;
    assign memory[  642 ] = 16'd27300;
    assign memory[  643 ] = 16'd27328;
    assign memory[  644 ] = 16'd27356;
    assign memory[  645 ] = 16'd27384;
    assign memory[  646 ] = 16'd27411;
    assign memory[  647 ] = 16'd27439;
    assign memory[  648 ] = 16'd27466;
    assign memory[  649 ] = 16'd27493;
    assign memory[  650 ] = 16'd27521;
    assign memory[  651 ] = 16'd27548;
    assign memory[  652 ] = 16'd27575;
    assign memory[  653 ] = 16'd27602;
    assign memory[  654 ] = 16'd27629;
    assign memory[  655 ] = 16'd27656;
    assign memory[  656 ] = 16'd27683;
    assign memory[  657 ] = 16'd27710;
    assign memory[  658 ] = 16'd27737;
    assign memory[  659 ] = 16'd27764;
    assign memory[  660 ] = 16'd27790;
    assign memory[  661 ] = 16'd27817;
    assign memory[  662 ] = 16'd27843;
    assign memory[  663 ] = 16'd27870;
    assign memory[  664 ] = 16'd27896;
    assign memory[  665 ] = 16'd27923;
    assign memory[  666 ] = 16'd27949;
    assign memory[  667 ] = 16'd27975;
    assign memory[  668 ] = 16'd28001;
    assign memory[  669 ] = 16'd28027;
    assign memory[  670 ] = 16'd28053;
    assign memory[  671 ] = 16'd28079;
    assign memory[  672 ] = 16'd28105;
    assign memory[  673 ] = 16'd28131;
    assign memory[  674 ] = 16'd28157;
    assign memory[  675 ] = 16'd28182;
    assign memory[  676 ] = 16'd28208;
    assign memory[  677 ] = 16'd28234;
    assign memory[  678 ] = 16'd28259;
    assign memory[  679 ] = 16'd28284;
    assign memory[  680 ] = 16'd28310;
    assign memory[  681 ] = 16'd28335;
    assign memory[  682 ] = 16'd28360;
    assign memory[  683 ] = 16'd28385;
    assign memory[  684 ] = 16'd28411;
    assign memory[  685 ] = 16'd28436;
    assign memory[  686 ] = 16'd28460;
    assign memory[  687 ] = 16'd28485;
    assign memory[  688 ] = 16'd28510;
    assign memory[  689 ] = 16'd28535;
    assign memory[  690 ] = 16'd28560;
    assign memory[  691 ] = 16'd28584;
    assign memory[  692 ] = 16'd28609;
    assign memory[  693 ] = 16'd28633;
    assign memory[  694 ] = 16'd28658;
    assign memory[  695 ] = 16'd28682;
    assign memory[  696 ] = 16'd28706;
    assign memory[  697 ] = 16'd28730;
    assign memory[  698 ] = 16'd28755;
    assign memory[  699 ] = 16'd28779;
    assign memory[  700 ] = 16'd28803;
    assign memory[  701 ] = 16'd28827;
    assign memory[  702 ] = 16'd28850;
    assign memory[  703 ] = 16'd28874;
    assign memory[  704 ] = 16'd28898;
    assign memory[  705 ] = 16'd28922;
    assign memory[  706 ] = 16'd28945;
    assign memory[  707 ] = 16'd28969;
    assign memory[  708 ] = 16'd28992;
    assign memory[  709 ] = 16'd29016;
    assign memory[  710 ] = 16'd29039;
    assign memory[  711 ] = 16'd29062;
    assign memory[  712 ] = 16'd29085;
    assign memory[  713 ] = 16'd29108;
    assign memory[  714 ] = 16'd29131;
    assign memory[  715 ] = 16'd29154;
    assign memory[  716 ] = 16'd29177;
    assign memory[  717 ] = 16'd29200;
    assign memory[  718 ] = 16'd29223;
    assign memory[  719 ] = 16'd29246;
    assign memory[  720 ] = 16'd29268;
    assign memory[  721 ] = 16'd29291;
    assign memory[  722 ] = 16'd29313;
    assign memory[  723 ] = 16'd29336;
    assign memory[  724 ] = 16'd29358;
    assign memory[  725 ] = 16'd29380;
    assign memory[  726 ] = 16'd29403;
    assign memory[  727 ] = 16'd29425;
    assign memory[  728 ] = 16'd29447;
    assign memory[  729 ] = 16'd29469;
    assign memory[  730 ] = 16'd29491;
    assign memory[  731 ] = 16'd29513;
    assign memory[  732 ] = 16'd29534;
    assign memory[  733 ] = 16'd29556;
    assign memory[  734 ] = 16'd29578;
    assign memory[  735 ] = 16'd29599;
    assign memory[  736 ] = 16'd29621;
    assign memory[  737 ] = 16'd29642;
    assign memory[  738 ] = 16'd29664;
    assign memory[  739 ] = 16'd29685;
    assign memory[  740 ] = 16'd29706;
    assign memory[  741 ] = 16'd29728;
    assign memory[  742 ] = 16'd29749;
    assign memory[  743 ] = 16'd29770;
    assign memory[  744 ] = 16'd29791;
    assign memory[  745 ] = 16'd29812;
    assign memory[  746 ] = 16'd29832;
    assign memory[  747 ] = 16'd29853;
    assign memory[  748 ] = 16'd29874;
    assign memory[  749 ] = 16'd29894;
    assign memory[  750 ] = 16'd29915;
    assign memory[  751 ] = 16'd29936;
    assign memory[  752 ] = 16'd29956;
    assign memory[  753 ] = 16'd29976;
    assign memory[  754 ] = 16'd29997;
    assign memory[  755 ] = 16'd30017;
    assign memory[  756 ] = 16'd30037;
    assign memory[  757 ] = 16'd30057;
    assign memory[  758 ] = 16'd30077;
    assign memory[  759 ] = 16'd30097;
    assign memory[  760 ] = 16'd30117;
    assign memory[  761 ] = 16'd30136;
    assign memory[  762 ] = 16'd30156;
    assign memory[  763 ] = 16'd30176;
    assign memory[  764 ] = 16'd30195;
    assign memory[  765 ] = 16'd30215;
    assign memory[  766 ] = 16'd30234;
    assign memory[  767 ] = 16'd30253;
    assign memory[  768 ] = 16'd30273;
    assign memory[  769 ] = 16'd30292;
    assign memory[  770 ] = 16'd30311;
    assign memory[  771 ] = 16'd30330;
    assign memory[  772 ] = 16'd30349;
    assign memory[  773 ] = 16'd30368;
    assign memory[  774 ] = 16'd30387;
    assign memory[  775 ] = 16'd30406;
    assign memory[  776 ] = 16'd30424;
    assign memory[  777 ] = 16'd30443;
    assign memory[  778 ] = 16'd30462;
    assign memory[  779 ] = 16'd30480;
    assign memory[  780 ] = 16'd30498;
    assign memory[  781 ] = 16'd30517;
    assign memory[  782 ] = 16'd30535;
    assign memory[  783 ] = 16'd30553;
    assign memory[  784 ] = 16'd30571;
    assign memory[  785 ] = 16'd30589;
    assign memory[  786 ] = 16'd30607;
    assign memory[  787 ] = 16'd30625;
    assign memory[  788 ] = 16'd30643;
    assign memory[  789 ] = 16'd30661;
    assign memory[  790 ] = 16'd30679;
    assign memory[  791 ] = 16'd30696;
    assign memory[  792 ] = 16'd30714;
    assign memory[  793 ] = 16'd30731;
    assign memory[  794 ] = 16'd30749;
    assign memory[  795 ] = 16'd30766;
    assign memory[  796 ] = 16'd30783;
    assign memory[  797 ] = 16'd30800;
    assign memory[  798 ] = 16'd30818;
    assign memory[  799 ] = 16'd30835;
    assign memory[  800 ] = 16'd30852;
    assign memory[  801 ] = 16'd30868;
    assign memory[  802 ] = 16'd30885;
    assign memory[  803 ] = 16'd30902;
    assign memory[  804 ] = 16'd30919;
    assign memory[  805 ] = 16'd30935;
    assign memory[  806 ] = 16'd30952;
    assign memory[  807 ] = 16'd30968;
    assign memory[  808 ] = 16'd30985;
    assign memory[  809 ] = 16'd31001;
    assign memory[  810 ] = 16'd31017;
    assign memory[  811 ] = 16'd31033;
    assign memory[  812 ] = 16'd31050;
    assign memory[  813 ] = 16'd31066;
    assign memory[  814 ] = 16'd31082;
    assign memory[  815 ] = 16'd31097;
    assign memory[  816 ] = 16'd31113;
    assign memory[  817 ] = 16'd31129;
    assign memory[  818 ] = 16'd31145;
    assign memory[  819 ] = 16'd31160;
    assign memory[  820 ] = 16'd31176;
    assign memory[  821 ] = 16'd31191;
    assign memory[  822 ] = 16'd31206;
    assign memory[  823 ] = 16'd31222;
    assign memory[  824 ] = 16'd31237;
    assign memory[  825 ] = 16'd31252;
    assign memory[  826 ] = 16'd31267;
    assign memory[  827 ] = 16'd31282;
    assign memory[  828 ] = 16'd31297;
    assign memory[  829 ] = 16'd31312;
    assign memory[  830 ] = 16'd31327;
    assign memory[  831 ] = 16'd31341;
    assign memory[  832 ] = 16'd31356;
    assign memory[  833 ] = 16'd31371;
    assign memory[  834 ] = 16'd31385;
    assign memory[  835 ] = 16'd31400;
    assign memory[  836 ] = 16'd31414;
    assign memory[  837 ] = 16'd31428;
    assign memory[  838 ] = 16'd31442;
    assign memory[  839 ] = 16'd31456;
    assign memory[  840 ] = 16'd31470;
    assign memory[  841 ] = 16'd31484;
    assign memory[  842 ] = 16'd31498;
    assign memory[  843 ] = 16'd31512;
    assign memory[  844 ] = 16'd31526;
    assign memory[  845 ] = 16'd31539;
    assign memory[  846 ] = 16'd31553;
    assign memory[  847 ] = 16'd31567;
    assign memory[  848 ] = 16'd31580;
    assign memory[  849 ] = 16'd31593;
    assign memory[  850 ] = 16'd31607;
    assign memory[  851 ] = 16'd31620;
    assign memory[  852 ] = 16'd31633;
    assign memory[  853 ] = 16'd31646;
    assign memory[  854 ] = 16'd31659;
    assign memory[  855 ] = 16'd31672;
    assign memory[  856 ] = 16'd31685;
    assign memory[  857 ] = 16'd31698;
    assign memory[  858 ] = 16'd31710;
    assign memory[  859 ] = 16'd31723;
    assign memory[  860 ] = 16'd31736;
    assign memory[  861 ] = 16'd31748;
    assign memory[  862 ] = 16'd31760;
    assign memory[  863 ] = 16'd31773;
    assign memory[  864 ] = 16'd31785;
    assign memory[  865 ] = 16'd31797;
    assign memory[  866 ] = 16'd31809;
    assign memory[  867 ] = 16'd31821;
    assign memory[  868 ] = 16'd31833;
    assign memory[  869 ] = 16'd31845;
    assign memory[  870 ] = 16'd31857;
    assign memory[  871 ] = 16'd31869;
    assign memory[  872 ] = 16'd31880;
    assign memory[  873 ] = 16'd31892;
    assign memory[  874 ] = 16'd31903;
    assign memory[  875 ] = 16'd31915;
    assign memory[  876 ] = 16'd31926;
    assign memory[  877 ] = 16'd31937;
    assign memory[  878 ] = 16'd31949;
    assign memory[  879 ] = 16'd31960;
    assign memory[  880 ] = 16'd31971;
    assign memory[  881 ] = 16'd31982;
    assign memory[  882 ] = 16'd31993;
    assign memory[  883 ] = 16'd32004;
    assign memory[  884 ] = 16'd32014;
    assign memory[  885 ] = 16'd32025;
    assign memory[  886 ] = 16'd32036;
    assign memory[  887 ] = 16'd32046;
    assign memory[  888 ] = 16'd32057;
    assign memory[  889 ] = 16'd32067;
    assign memory[  890 ] = 16'd32077;
    assign memory[  891 ] = 16'd32087;
    assign memory[  892 ] = 16'd32098;
    assign memory[  893 ] = 16'd32108;
    assign memory[  894 ] = 16'd32118;
    assign memory[  895 ] = 16'd32128;
    assign memory[  896 ] = 16'd32137;
    assign memory[  897 ] = 16'd32147;
    assign memory[  898 ] = 16'd32157;
    assign memory[  899 ] = 16'd32166;
    assign memory[  900 ] = 16'd32176;
    assign memory[  901 ] = 16'd32185;
    assign memory[  902 ] = 16'd32195;
    assign memory[  903 ] = 16'd32204;
    assign memory[  904 ] = 16'd32213;
    assign memory[  905 ] = 16'd32223;
    assign memory[  906 ] = 16'd32232;
    assign memory[  907 ] = 16'd32241;
    assign memory[  908 ] = 16'd32250;
    assign memory[  909 ] = 16'd32258;
    assign memory[  910 ] = 16'd32267;
    assign memory[  911 ] = 16'd32276;
    assign memory[  912 ] = 16'd32285;
    assign memory[  913 ] = 16'd32293;
    assign memory[  914 ] = 16'd32302;
    assign memory[  915 ] = 16'd32310;
    assign memory[  916 ] = 16'd32318;
    assign memory[  917 ] = 16'd32327;
    assign memory[  918 ] = 16'd32335;
    assign memory[  919 ] = 16'd32343;
    assign memory[  920 ] = 16'd32351;
    assign memory[  921 ] = 16'd32359;
    assign memory[  922 ] = 16'd32367;
    assign memory[  923 ] = 16'd32375;
    assign memory[  924 ] = 16'd32382;
    assign memory[  925 ] = 16'd32390;
    assign memory[  926 ] = 16'd32397;
    assign memory[  927 ] = 16'd32405;
    assign memory[  928 ] = 16'd32412;
    assign memory[  929 ] = 16'd32420;
    assign memory[  930 ] = 16'd32427;
    assign memory[  931 ] = 16'd32434;
    assign memory[  932 ] = 16'd32441;
    assign memory[  933 ] = 16'd32448;
    assign memory[  934 ] = 16'd32455;
    assign memory[  935 ] = 16'd32462;
    assign memory[  936 ] = 16'd32469;
    assign memory[  937 ] = 16'd32476;
    assign memory[  938 ] = 16'd32482;
    assign memory[  939 ] = 16'd32489;
    assign memory[  940 ] = 16'd32495;
    assign memory[  941 ] = 16'd32502;
    assign memory[  942 ] = 16'd32508;
    assign memory[  943 ] = 16'd32514;
    assign memory[  944 ] = 16'd32521;
    assign memory[  945 ] = 16'd32527;
    assign memory[  946 ] = 16'd32533;
    assign memory[  947 ] = 16'd32539;
    assign memory[  948 ] = 16'd32545;
    assign memory[  949 ] = 16'd32550;
    assign memory[  950 ] = 16'd32556;
    assign memory[  951 ] = 16'd32562;
    assign memory[  952 ] = 16'd32567;
    assign memory[  953 ] = 16'd32573;
    assign memory[  954 ] = 16'd32578;
    assign memory[  955 ] = 16'd32584;
    assign memory[  956 ] = 16'd32589;
    assign memory[  957 ] = 16'd32594;
    assign memory[  958 ] = 16'd32599;
    assign memory[  959 ] = 16'd32604;
    assign memory[  960 ] = 16'd32609;
    assign memory[  961 ] = 16'd32614;
    assign memory[  962 ] = 16'd32619;
    assign memory[  963 ] = 16'd32624;
    assign memory[  964 ] = 16'd32628;
    assign memory[  965 ] = 16'd32633;
    assign memory[  966 ] = 16'd32637;
    assign memory[  967 ] = 16'd32642;
    assign memory[  968 ] = 16'd32646;
    assign memory[  969 ] = 16'd32650;
    assign memory[  970 ] = 16'd32655;
    assign memory[  971 ] = 16'd32659;
    assign memory[  972 ] = 16'd32663;
    assign memory[  973 ] = 16'd32667;
    assign memory[  974 ] = 16'd32671;
    assign memory[  975 ] = 16'd32674;
    assign memory[  976 ] = 16'd32678;
    assign memory[  977 ] = 16'd32682;
    assign memory[  978 ] = 16'd32685;
    assign memory[  979 ] = 16'd32689;
    assign memory[  980 ] = 16'd32692;
    assign memory[  981 ] = 16'd32696;
    assign memory[  982 ] = 16'd32699;
    assign memory[  983 ] = 16'd32702;
    assign memory[  984 ] = 16'd32705;
    assign memory[  985 ] = 16'd32708;
    assign memory[  986 ] = 16'd32711;
    assign memory[  987 ] = 16'd32714;
    assign memory[  988 ] = 16'd32717;
    assign memory[  989 ] = 16'd32720;
    assign memory[  990 ] = 16'd32722;
    assign memory[  991 ] = 16'd32725;
    assign memory[  992 ] = 16'd32728;
    assign memory[  993 ] = 16'd32730;
    assign memory[  994 ] = 16'd32732;
    assign memory[  995 ] = 16'd32735;
    assign memory[  996 ] = 16'd32737;
    assign memory[  997 ] = 16'd32739;
    assign memory[  998 ] = 16'd32741;
    assign memory[  999 ] = 16'd32743;
    assign memory[ 1000 ] = 16'd32745;
    assign memory[ 1001 ] = 16'd32747;
    assign memory[ 1002 ] = 16'd32748;
    assign memory[ 1003 ] = 16'd32750;
    assign memory[ 1004 ] = 16'd32752;
    assign memory[ 1005 ] = 16'd32753;
    assign memory[ 1006 ] = 16'd32755;
    assign memory[ 1007 ] = 16'd32756;
    assign memory[ 1008 ] = 16'd32757;
    assign memory[ 1009 ] = 16'd32758;
    assign memory[ 1010 ] = 16'd32759;
    assign memory[ 1011 ] = 16'd32760;
    assign memory[ 1012 ] = 16'd32761;
    assign memory[ 1013 ] = 16'd32762;
    assign memory[ 1014 ] = 16'd32763;
    assign memory[ 1015 ] = 16'd32764;
    assign memory[ 1016 ] = 16'd32765;
    assign memory[ 1017 ] = 16'd32765;
    assign memory[ 1018 ] = 16'd32766;
    assign memory[ 1019 ] = 16'd32766;
    assign memory[ 1020 ] = 16'd32766;
    assign memory[ 1021 ] = 16'd32767;
    assign memory[ 1022 ] = 16'd32767;
    assign memory[ 1023 ] = 16'd32767;

endmodule
