
module note_address (
	input 		[5:0] 	note,
	output reg	[44:0] 	note_addr
);
	always @(note)
		case (note) // 1:octave 2:note 3:sharp 4:note 5:flat *32 is blank space
			6'd00: note_addr = {(9'd18 << 3), (9'd05 << 3), (9'd19 << 3), (9'd20 << 3), (9'd32 << 3)}; // REST
			6'd01: note_addr = {(9'd49 << 3), (9'd01 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 1A
			6'd02: note_addr = {(9'd49 << 3), (9'd01 << 3), (9'd35 << 3), (9'd02 << 3), (9'd63 << 3)}; // 1A#Bb
			6'd03: note_addr = {(9'd49 << 3), (9'd02 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 1B
			6'd04: note_addr = {(9'd49 << 3), (9'd03 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 1C
			6'd05: note_addr = {(9'd49 << 3), (9'd03 << 3), (9'd35 << 3), (9'd04 << 3), (9'd63 << 3)}; // 1C#Db
			6'd06: note_addr = {(9'd49 << 3), (9'd04 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 1D
			6'd07: note_addr = {(9'd49 << 3), (9'd04 << 3), (9'd35 << 3), (9'd05 << 3), (9'd63 << 3)}; // 1D#Eb
			6'd08: note_addr = {(9'd49 << 3), (9'd05 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 1E
			6'd09: note_addr = {(9'd49 << 3), (9'd06 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 1F
			6'd10: note_addr = {(9'd49 << 3), (9'd06 << 3), (9'd35 << 3), (9'd07 << 3), (9'd63 << 3)}; // 1F#Gb
			6'd11: note_addr = {(9'd49 << 3), (9'd07 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 1G
			6'd12: note_addr = {(9'd49 << 3), (9'd07 << 3), (9'd35 << 3), (9'd01 << 3), (9'd63 << 3)}; // 1G#Ab
			6'd13: note_addr = {(9'd50 << 3), (9'd01 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 2A
			6'd14: note_addr = {(9'd50 << 3), (9'd01 << 3), (9'd35 << 3), (9'd02 << 3), (9'd63 << 3)}; // 2A#Bb
			6'd15: note_addr = {(9'd50 << 3), (9'd02 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 2B
			6'd16: note_addr = {(9'd50 << 3), (9'd03 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 2C
			6'd17: note_addr = {(9'd50 << 3), (9'd03 << 3), (9'd35 << 3), (9'd04 << 3), (9'd63 << 3)}; // 2C#Db
			6'd18: note_addr = {(9'd50 << 3), (9'd04 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 2D
			6'd19: note_addr = {(9'd50 << 3), (9'd04 << 3), (9'd35 << 3), (9'd05 << 3), (9'd63 << 3)}; // 2D#Eb
			6'd20: note_addr = {(9'd50 << 3), (9'd05 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 2E
			6'd21: note_addr = {(9'd50 << 3), (9'd06 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 2F
			6'd22: note_addr = {(9'd50 << 3), (9'd06 << 3), (9'd35 << 3), (9'd07 << 3), (9'd63 << 3)}; // 2F#Gb
			6'd23: note_addr = {(9'd50 << 3), (9'd07 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 2G
			6'd24: note_addr = {(9'd50 << 3), (9'd07 << 3), (9'd35 << 3), (9'd01 << 3), (9'd63 << 3)}; // 2G#Ab
			6'd25: note_addr = {(9'd51 << 3), (9'd01 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 3A
			6'd26: note_addr = {(9'd51 << 3), (9'd01 << 3), (9'd35 << 3), (9'd02 << 3), (9'd63 << 3)}; // 3A#Bb
			6'd27: note_addr = {(9'd51 << 3), (9'd02 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 3B
			6'd63: note_addr = {(9'd51 << 3), (9'd03 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 3C
			6'd29: note_addr = {(9'd51 << 3), (9'd03 << 3), (9'd35 << 3), (9'd04 << 3), (9'd63 << 3)}; // 3C#Db
			6'd30: note_addr = {(9'd51 << 3), (9'd04 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 3D
			6'd31: note_addr = {(9'd51 << 3), (9'd04 << 3), (9'd35 << 3), (9'd05 << 3), (9'd63 << 3)}; // 3D#Eb
			6'd32: note_addr = {(9'd51 << 3), (9'd05 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 3E
			6'd33: note_addr = {(9'd51 << 3), (9'd06 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 3F
			6'd34: note_addr = {(9'd51 << 3), (9'd06 << 3), (9'd35 << 3), (9'd07 << 3), (9'd63 << 3)}; // 3F#Gb
			6'd35: note_addr = {(9'd51 << 3), (9'd07 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 3G
			6'd36: note_addr = {(9'd51 << 3), (9'd07 << 3), (9'd35 << 3), (9'd01 << 3), (9'd63 << 3)}; // 3G#Ab
			6'd37: note_addr = {(9'd52 << 3), (9'd01 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 4A
			6'd38: note_addr = {(9'd52 << 3), (9'd01 << 3), (9'd35 << 3), (9'd02 << 3), (9'd63 << 3)}; // 4A#Bb
			6'd39: note_addr = {(9'd52 << 3), (9'd02 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 4B
			6'd40: note_addr = {(9'd52 << 3), (9'd03 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 4C
			6'd41: note_addr = {(9'd52 << 3), (9'd03 << 3), (9'd35 << 3), (9'd04 << 3), (9'd63 << 3)}; // 4C#Db
			6'd42: note_addr = {(9'd52 << 3), (9'd04 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 4D
			6'd43: note_addr = {(9'd52 << 3), (9'd04 << 3), (9'd35 << 3), (9'd05 << 3), (9'd63 << 3)}; // 4D#Eb
			6'd44: note_addr = {(9'd52 << 3), (9'd05 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 4E
			6'd45: note_addr = {(9'd52 << 3), (9'd06 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 4F
			6'd46: note_addr = {(9'd52 << 3), (9'd06 << 3), (9'd35 << 3), (9'd07 << 3), (9'd63 << 3)}; // 4F#Gb
			6'd47: note_addr = {(9'd52 << 3), (9'd07 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 4G
			6'd48: note_addr = {(9'd52 << 3), (9'd07 << 3), (9'd35 << 3), (9'd01 << 3), (9'd63 << 3)}; // 4G#Ab
			6'd49: note_addr = {(9'd53 << 3), (9'd01 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 5A
			6'd50: note_addr = {(9'd53 << 3), (9'd01 << 3), (9'd35 << 3), (9'd02 << 3), (9'd63 << 3)}; // 5A#Bb
			6'd51: note_addr = {(9'd53 << 3), (9'd02 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 5B
			6'd52: note_addr = {(9'd53 << 3), (9'd03 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 5C
			6'd53: note_addr = {(9'd53 << 3), (9'd03 << 3), (9'd35 << 3), (9'd04 << 3), (9'd63 << 3)}; // 5C#Db
			6'd54: note_addr = {(9'd53 << 3), (9'd04 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 5D
			6'd55: note_addr = {(9'd53 << 3), (9'd04 << 3), (9'd35 << 3), (9'd05 << 3), (9'd63 << 3)}; // 5D#Eb
			6'd56: note_addr = {(9'd53 << 3), (9'd05 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 5E
			6'd57: note_addr = {(9'd53 << 3), (9'd06 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 5F
			6'd58: note_addr = {(9'd53 << 3), (9'd06 << 3), (9'd35 << 3), (9'd07 << 3), (9'd63 << 3)}; // 5F#Gb
			6'd59: note_addr = {(9'd53 << 3), (9'd07 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 5G
			6'd60: note_addr = {(9'd53 << 3), (9'd07 << 3), (9'd35 << 3), (9'd01 << 3), (9'd63 << 3)}; // 5G#Ab
			6'd61: note_addr = {(9'd54 << 3), (9'd01 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 6A
			6'd62: note_addr = {(9'd54 << 3), (9'd01 << 3), (9'd35 << 3), (9'd02 << 3), (9'd63 << 3)}; // 6A#Bb
			6'd63: note_addr = {(9'd54 << 3), (9'd02 << 3), (9'd32 << 3), (9'd32 << 3), (9'd32 << 3)}; // 6B
			default: note_addr = {5{(9'd32 << 3)}};
		endcase
		
endmodule
